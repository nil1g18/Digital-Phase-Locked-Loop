`define N_BIT 16